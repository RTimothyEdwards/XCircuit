**********
LZ_0 1 int_node0_2 int_node1_1 1.2121
