************
RZ_0 1 2 1.92517e-11
