* standard_cells.cir, netlists for verifying standard cells
* Conrad Ziesler and Tim Edwards, MultiGiG, Inc.
* Standard cells are from the IIT standard cell library.

.subckt MUX2X1 vdd gnd A B Y S
M1 x1 A gnd gnd nfet l=180n w=1.80u m=1
M2 x2 A vdd vdd pfet l=180n w=3.60u m=1
M3 x2 S Y vdd pfet l=180n w=3.60u m=1
M4 x1 sbar Y gnd nfet l=180n w=1.80u m=1
M5 sbar S vdd vdd pfet l=180n w=1.80u m=1
M6 sbar S gnd gnd nfet l=180n w=0.90u m=1
M7 Y sbar x3 vdd pfet l=180n w=3.60u m=1
M8 Y S x4 gnd nfet l=180n w=1.80u m=1
M9 x3 B vdd vdd pfet l=180n w=3.60u m=1
M10 x4 B gnd gnd nfet l=180n w=1.80u m=1
.ends

.subckt TBUFX2 vdd gnd A Y En
M1 enb En gnd gnd nfet l=180n w=1.80u m=1
M2 enb En vdd vdd pfet l=180n w=3.60u m=1
M4 i A vdd vdd pfet l=180n w=3.60u m=2
M3 i enb Y vdd pfet l=180n w=3.60u m=2
M5 j En Y gnd nfet l=180n w=1.80u m=2
M6 j A gnd gnd nfet l=180n w=1.80u m=2
.ends

.subckt BUFX4 vdd gnd A Y
M1 x A gnd gnd nfet l=180n w=1.35u m=1
M2 x A vdd vdd pfet l=180n w=2.70u m=1
M3 Y x gnd gnd nfet l=180n w=1.80u m=2
M4 Y x vdd vdd pfet l=180n w=3.60u m=2
.ends

.subckt BUFX2 vdd gnd A Y
M1 x A gnd gnd nfet l=180n w=0.90u m=1
M2 x A vdd vdd pfet l=180n w=1.80u m=1
M3 Y x gnd gnd nfet l=180n w=1.80u m=1
M4 Y x vdd vdd pfet l=180n w=3.60u m=1
.ends

.subckt INVX1 vdd gnd A Y
M1 Y A gnd gnd nfet l=180n w=0.90u m=1
M2 Y A vdd vdd pfet l=180n w=1.80u m=1
.ends

.subckt INVX2 vdd gnd A Y
M1 Y A gnd gnd nfet l=180n w=1.80u m=1
M2 Y A vdd vdd pfet l=180n w=3.60u m=1
.ends

.subckt NOR2X1 vdd gnd A B Y
M1 Y A gnd gnd nfet l=180n w=0.90u m=1
M2 Y B gnd gnd nfet l=180n w=0.90u m=1
M3 x1 A vdd vdd pfet l=180n w=3.60u m=1
M4 Y  B x1  vdd pfet l=180n w=3.60u m=1
.ends

.subckt NOR3X1 vdd gnd A B C Y
M1 Y A gnd gnd nfet l=180n w=0.90u m=1
M2 Y B gnd gnd nfet l=180n w=0.90u m=1
M3 Y C gnd gnd nfet l=180n w=0.90u m=1
M4 x1 A vdd vdd pfet l=180n w=2.70u m=2
M5 x2 B x1  vdd pfet l=180n w=2.70u m=2
M6 Y  C x2  vdd pfet l=180n w=2.70u m=2
.ends

.subckt NAND2X1 vdd gnd A B Y
M1 x1 A gnd gnd nfet l=180n w=1.80u m=1
M2 Y  B x1  gnd nfet l=180n w=1.80u m=1
M3 Y  A vdd vdd pfet l=180n w=1.80u m=1
M4 Y  B vdd vdd pfet l=180n w=1.80u m=1
.ends

.subckt NAND3X1 vdd gnd A B C Y
M1 x1 A gnd gnd nfet l=180n w=2.70u m=1
M2 x2 B x1  gnd nfet l=180n w=2.70u m=1
M3 Y  C x2  gnd nfet l=180n w=2.70u m=1
M4 Y  A vdd vdd pfet l=180n w=1.80u m=1
M5 Y  B vdd vdd pfet l=180n w=1.80u m=1
M6 Y  C vdd vdd pfet l=180n w=1.80u m=1
.ends

.subckt OR2X1 vdd gnd A B Y
M1 x2 A gnd gnd nfet l=180n w=0.90u m=1
M2 x2 B gnd gnd nfet l=180n w=0.90u m=1
M3 x1 B vdd vdd pfet l=180n w=3.60u m=1
M4 x2 A x1  vdd pfet l=180n w=3.60u m=1
M5 Y x2 gnd gnd nfet l=180n w=0.90u m=1
M6 Y x2 vdd vdd pfet l=180n w=1.80u m=1
.ends

.subckt LATCH vdd gnd CLK D Q
M1 cb CLK gnd gnd nfet l=180n w=0.90u m=2
M2 cb CLK vdd vdd pfet l=180n w=0.90u m=4

M3 x2 D  vdd vdd pfet l=180n w=0.90u m=2
M4 qb cb   x2  vdd pfet l=180n w=0.90u m=2
M5 x4 D  gnd  gnd nfet l=180n w=0.90u m=1
M6 qb CLK   x4   gnd nfet l=180n w=0.90u m=1

M7  x5 Q  vdd vdd pfet l=180n w=0.90u m=1
M8  qb CLK    x5  vdd pfet l=180n w=0.90u m=1
M9  x7 Q   gnd  gnd nfet l=180n w=0.90u m=1
M10 qb cb    x7   gnd nfet l=180n w=0.90u m=1

M11 Q qb gnd gnd nfet l=180n w=0.90u m=2
M12 Q qb vdd vdd pfet l=180n w=0.90u m=4
.ends
