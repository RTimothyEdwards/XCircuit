* LZ_0 1 int_node0_2 1.92517e-11
.END
